library ieee;
use ieee.std_logic_1164.all;

entity eq is
	port(
		eq1: in std_logic_vector(15 downto 0);
		eq2: in std_logic_vector(15 downto 0);
		eq_out: out std_logic)
end entity;

architecture arch of eq is
begin
	
	eq_out <= '1' when eq_1 = eq_2 else '0';

end architecture;